//------Lab2 Comparator
module comparator(
    input [3:0] V,
    output z
);
    assign z = V[3];
endmodule